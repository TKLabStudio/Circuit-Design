library verilog;
use verilog.vl_types.all;
entity P1041217_vlg_vec_tst is
end P1041217_vlg_vec_tst;
