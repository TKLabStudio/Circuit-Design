library verilog;
use verilog.vl_types.all;
entity P1041217 is
    port(
        o0              : out    vl_logic;
        CLK             : in     vl_logic;
        BUTT            : in     vl_logic;
        o1              : out    vl_logic;
        o2              : out    vl_logic;
        o3              : out    vl_logic;
        o4              : out    vl_logic;
        o5              : out    vl_logic;
        o6              : out    vl_logic;
        o7              : out    vl_logic;
        o8              : out    vl_logic;
        o9              : out    vl_logic
    );
end P1041217;
